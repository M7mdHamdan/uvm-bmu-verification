class BmuSequencer extends uvm_sequencer;
    `uvm_utils_

    function new (string name = "BmuSequencer");
        super.new(name);
    endfunction;


endclass: BmuSequencer