`define RV_INST_ACCESS_MASK5 'hffffffff
`define RV_DATA_ACCESS_ENABLE4 1'h0
`define RV_INST_ACCESS_ENABLE3 1'h0
`define RV_INST_ACCESS_ENABLE0 1'h0
`define RV_INST_ACCESS_MASK3 'hffffffff
`define RV_DATA_ACCESS_ENABLE5 1'h0
`define RV_DATA_ACCESS_MASK5 'hffffffff
`define RV_DATA_ACCESS_ADDR3 'h00000000
`define RV_INST_ACCESS_ENABLE7 1'h0
`define RV_DATA_ACCESS_ADDR6 'h00000000
`define RV_INST_ACCESS_MASK7 'hffffffff
`define RV_INST_ACCESS_ENABLE6 1'h0
`define RV_INST_ACCESS_ENABLE5 1'h0
`define RV_DATA_ACCESS_ADDR4 'h00000000
`define RV_DATA_ACCESS_ADDR7 'h00000000
`define RV_DATA_ACCESS_MASK3 'hffffffff
`define RV_INST_ACCESS_MASK4 'hffffffff
`define RV_DATA_ACCESS_ADDR1 'h00000000
`define RV_INST_ACCESS_ADDR4 'h00000000
`define RV_INST_ACCESS_ADDR3 'h00000000
`define RV_DATA_ACCESS_ENABLE1 1'h0
`define RV_DATA_ACCESS_ADDR0 'h00000000
`define RV_DATA_ACCESS_MASK0 'hffffffff
`define RV_DATA_ACCESS_MASK6 'hffffffff
`define RV_INST_ACCESS_ADDR7 'h00000000
`define RV_INST_ACCESS_MASK0 'hffffffff
`define RV_DATA_ACCESS_ADDR5 'h00000000
`define RV_DATA_ACCESS_ADDR2 'h00000000
`define RV_DATA_ACCESS_MASK4 'hffffffff
`define RV_DATA_ACCESS_MASK1 'hffffffff
`define RV_INST_ACCESS_ADDR0 'h00000000
`define RV_INST_ACCESS_ADDR2 'h00000000
`define RV_DATA_ACCESS_ENABLE0 1'h0
`define RV_DATA_ACCESS_ENABLE2 1'h0
`define RV_DATA_ACCESS_ENABLE7 1'h0
`define RV_INST_ACCESS_ENABLE4 1'h0
`define RV_DATA_ACCESS_MASK7 'hffffffff
`define RV_INST_ACCESS_ADDR5 'h00000000
`define RV_DATA_ACCESS_MASK2 'hffffffff
`define RV_INST_ACCESS_ENABLE1 1'h0
`define RV_INST_ACCESS_MASK6 'hffffffff
`define RV_DATA_ACCESS_ENABLE3 1'h0
`define RV_INST_ACCESS_ADDR6 'h00000000
`define RV_INST_ACCESS_MASK2 'hffffffff
`define RV_INST_ACCESS_ENABLE2 1'h0
`define RV_DATA_ACCESS_ENABLE6 1'h0
`define RV_INST_ACCESS_ADDR1 'h00000000
`define RV_INST_ACCESS_MASK1 'hffffffff
`define RV_LSU2DMA 0
`define RV_BITMANIP_ZBR 0
`define RV_BITMANIP_ZBP 0
`define RV_BITMANIP_ZBF 0
`define RV_BITMANIP_ZBC 1
`define RV_BITMANIP_ZBA 1
`define RV_DIV_NEW 1
`define RV_BITMANIP_ZBE 0
`define RV_DIV_BIT 4
`define RV_LSU_NUM_NBLOAD 4
`define RV_BITMANIP_ZBB 1
`define RV_FPGA_OPTIMIZE 1
`define RV_BITMANIP_ZBS 1
`define RV_FAST_INTERRUPT_REDIRECT 1
`define RV_DMA_BUF_DEPTH 5
`define RV_LSU_STBUF_DEPTH 4
`define RV_LSU_NUM_NBLOAD_WIDTH 2
`define RV_TIMER_LEGAL_EN 1
`define RV_ICCM_ICACHE 1
`define RV_IFU_BUS_TAG 3
`define RV_LSU_BUS_ID 1
`define RV_LSU_BUS_TAG 3
`define RV_SB_BUS_ID 1
`define RV_DMA_BUS_ID 1
`define RV_IFU_BUS_PRTY 2
`define RV_SB_BUS_PRTY 2
`define RV_LSU_BUS_PRTY 2
`define RV_SB_BUS_TAG 1
`define RV_IFU_BUS_ID 1
`define RV_DMA_BUS_PRTY 2
`define RV_BUS_PRTY_DEFAULT 2'h3
`define RV_DMA_BUS_TAG 1
`define RV_DCCM_WIDTH_BITS 2
`define RV_DCCM_REGION 4'hf
`define RV_DCCM_RESERVED 'h1400
`define RV_DCCM_SIZE 64
`define RV_DCCM_DATA_WIDTH 32
`define RV_DCCM_FDATA_WIDTH 39
`define RV_DCCM_BYTE_WIDTH 4
`define RV_DCCM_DATA_CELL ram_4096x39
`define RV_DCCM_ENABLE 1
`define RV_DCCM_BITS 16
`define RV_DCCM_OFFSET 28'h40000
`define RV_DCCM_ECC_WIDTH 7
`define RV_DCCM_SIZE_64 
`define RV_DCCM_ROWS 4096
`define RV_DCCM_BANK_BITS 2
`define RV_DCCM_NUM_BANKS 4
`define RV_DCCM_INDEX_BITS 12
`define RV_LSU_SB_BITS 16
`define RV_DCCM_EADR 32'hf004ffff
`define RV_DCCM_NUM_BANKS_4 
`define RV_DCCM_SADR 32'hf0040000
`define RV_RESET_VEC 'h80000000
`define RV_RET_STACK_SIZE 8
`define RV_XLEN 32
`define RV_TARGET default
`define RV_BTB_BTAG_FOLD 0
`define RV_BTB_INDEX3_HI 25
`define RV_BTB_INDEX3_LO 18
`define RV_BTB_INDEX1_LO 2
`define RV_BTB_ENABLE 1
`define RV_BTB_ADDR_HI 9
`define RV_BTB_FOLD2_INDEX_HASH 0
`define RV_BTB_INDEX2_HI 17
`define RV_BTB_INDEX1_HI 9
`define RV_BTB_ADDR_LO 2
`define RV_BTB_INDEX2_LO 10
`define RV_BTB_ARRAY_DEPTH 256
`define RV_BTB_BTAG_SIZE 5
`define RV_BTB_SIZE 512
`define RV_BTB_TOFFSET_SIZE 12
`define RV_ICCM_BANK_HI 3
`define RV_ICCM_ENABLE 1
`define RV_ICCM_BITS 16
`define RV_ICCM_OFFSET 10'he000000
`define RV_ICCM_SADR 32'hee000000
`define RV_ICCM_DATA_CELL ram_4096x39
`define RV_ICCM_NUM_BANKS_4 
`define RV_ICCM_EADR 32'hee00ffff
`define RV_ICCM_BANK_INDEX_LO 4
`define RV_ICCM_NUM_BANKS 4
`define RV_ICCM_BANK_BITS 2
`define RV_ICCM_ROWS 4096
`define RV_ICCM_REGION 4'he
`define RV_ICCM_RESERVED 'h1000
`define RV_ICCM_SIZE_64 
`define RV_ICCM_INDEX_BITS 12
`define RV_ICCM_SIZE 64
`define RV_ICACHE_TAG_INDEX_LO 6
`define RV_ICACHE_DATA_DEPTH 512
`define RV_ICACHE_SCND_LAST 6
`define RV_ICACHE_ECC 1
`define RV_ICACHE_TAG_NUM_BYPASS_WIDTH 2
`define RV_ICACHE_DATA_WIDTH 64
`define RV_ICACHE_BEAT_ADDR_HI 5
`define RV_ICACHE_NUM_WAYS 2
`define RV_ICACHE_BYPASS_ENABLE 1
`define RV_ICACHE_WAYPACK 1
`define RV_ICACHE_INDEX_HI 12
`define RV_ICACHE_BANKS_WAY 2
`define RV_ICACHE_SIZE 16
`define RV_ICACHE_TAG_BYPASS_ENABLE 1
`define RV_ICACHE_NUM_BYPASS 2
`define RV_ICACHE_TAG_CELL ram_128x25
`define RV_ICACHE_TAG_DEPTH 128
`define RV_ICACHE_BANK_WIDTH 8
`define RV_ICACHE_BANK_LO 3
`define RV_ICACHE_NUM_LINES 256
`define RV_ICACHE_NUM_BEATS 8
`define RV_ICACHE_NUM_LINES_WAY 128
`define RV_ICACHE_TAG_LO 13
`define RV_ICACHE_BANK_HI 3
`define RV_ICACHE_ENABLE 1
`define RV_ICACHE_DATA_CELL ram_512x71
`define RV_ICACHE_NUM_LINES_BANK 64
`define RV_ICACHE_FDATA_WIDTH 71
`define RV_ICACHE_BEAT_BITS 3
`define RV_ICACHE_2BANKS 1
`define RV_ICACHE_TAG_NUM_BYPASS 2
`define RV_ICACHE_NUM_BYPASS_WIDTH 2
`define RV_ICACHE_STATUS_BITS 1
`define RV_ICACHE_BANK_BITS 1
`define RV_ICACHE_DATA_INDEX_LO 4
`define RV_ICACHE_LN_SZ 64
`define RV_UNUSED_REGION7 'h10000000
`define RV_UNUSED_REGION4 'h40000000
`define RV_UNUSED_REGION8 'h00000000
`define RV_SERIALIO 'hd0580000
`define RV_UNUSED_REGION2 'h60000000
`define RV_UNUSED_REGION1 'h70000000
`define RV_UNUSED_REGION0 'h90000000
`define RV_UNUSED_REGION3 'h50000000
`define RV_UNUSED_REGION5 'h30000000
`define RV_EXTERNAL_DATA_1 'hb0000000
`define RV_DEBUG_SB_MEM 'ha0580000
`define RV_UNUSED_REGION6 'h20000000
`define RV_EXTERNAL_DATA 'hc0580000
`define RV_NMI_VEC 'h11110000
`define RV_BHT_HASH_STRING {hashin[8+1:2]^ghr[8-1:0]}// cf2
`define RV_BHT_ADDR_HI 9
`define RV_BHT_GHR_RANGE 7:0
`define RV_BHT_GHR_HASH_1 
`define RV_BHT_GHR_SIZE 8
`define RV_BHT_SIZE 512
`define RV_BHT_ADDR_LO 2
`define RV_BHT_ARRAY_DEPTH 256
`define RV_NUMIREGS 32
`define RV_PIC_MEIPL_MASK 'hf
`define RV_PIC_MEIP_COUNT 1
`define RV_PIC_BITS 15
`define RV_PIC_REGION 4'hf
`define RV_PIC_INT_WORDS 1
`define RV_PIC_MEIE_COUNT 31
`define RV_PIC_MPICCFG_MASK 'h1
`define RV_PIC_TOTAL_INT_PLUS1 32
`define RV_PIC_MEIGWCTRL_MASK 'h3
`define RV_PIC_MEIP_OFFSET 'h1000
`define RV_PIC_BASE_ADDR 32'hf00c0000
`define RV_PIC_MEIPT_MASK 'h0
`define RV_PIC_MEIGWCTRL_OFFSET 'h4000
`define RV_PIC_MEIPL_OFFSET 'h0000
`define RV_PIC_MEIPT_COUNT 31
`define RV_PIC_TOTAL_INT 31
`define RV_PIC_MEIGWCLR_COUNT 31
`define RV_PIC_MPICCFG_COUNT 1
`define RV_PIC_SIZE 32
`define RV_PIC_MEIGWCTRL_COUNT 31
`define RV_PIC_MEIE_OFFSET 'h2000
`define RV_PIC_MEIPL_COUNT 31
`define RV_PIC_OFFSET 10'hc0000
`define RV_PIC_MEIP_MASK 'h0
`define RV_PIC_MEIPT_OFFSET 'h3004
`define RV_PIC_MEIGWCLR_MASK 'h0
`define RV_PIC_MEIE_MASK 'h1
`define RV_PIC_MPICCFG_OFFSET 'h3000
`define RV_PIC_MEIGWCLR_OFFSET 'h5000
`define RV_CONFIG_KEY 32'hdeadbeef
`define CLOCK_PERIOD 100
`define CPU_TOP `RV_TOP.orv
`define TOP tb_top
`define RV_BUILD_AXI4 1
`define RV_TOP `TOP.rvtop
`define RV_STERR_ROLLBACK 0
`define RV_EXT_ADDRWIDTH 32
`define RV_EXT_DATAWIDTH 64
`define SDVT_AHB 0
`define RV_LDERR_ROLLBACK 1
`define RV_ASSERT_ON 
`define RV_BUILD_AXI_NATIVE 1
`define TEC_RV_ICG clockhdr
`define REGWIDTH 32
parameter rtl_param_t pt = '{
	BHT_ADDR_HI            : 8'h09         ,
	BHT_ADDR_LO            : 6'h02         ,
	BHT_ARRAY_DEPTH        : 15'h0100       ,
	BHT_GHR_HASH_1         : 5'h00         ,
	BHT_GHR_SIZE           : 8'h08         ,
	BHT_SIZE               : 16'h0200       ,
	BITMANIP_ZBA           : 5'h01         ,
	BITMANIP_ZBB           : 5'h01         ,
	BITMANIP_ZBC           : 5'h01         ,
	BITMANIP_ZBE           : 5'h00         ,
	BITMANIP_ZBF           : 5'h00         , 
	BITMANIP_ZBP           : 5'h00         ,
	BITMANIP_ZBR           : 5'h00         ,
	BITMANIP_ZBS           : 5'h01         ,
	BTB_ADDR_HI            : 9'h009        ,
	BTB_ADDR_LO            : 6'h02         ,
	BTB_ARRAY_DEPTH        : 13'h0100      ,
	BTB_BTAG_FOLD          : 5'h00         ,
	BTB_BTAG_SIZE          : 9'h005        ,
	BTB_ENABLE             : 5'h01         ,
	BTB_FOLD2_INDEX_HASH   : 5'h00         ,
	BTB_FULLYA             : 5'h00         ,
	BTB_INDEX1_HI          : 9'h009        ,
	BTB_INDEX1_LO          : 9'h002        ,
	BTB_INDEX2_HI          : 9'h011        ,
	BTB_INDEX2_LO          : 9'h00A        ,
	BTB_INDEX3_HI          : 9'h019        ,
	BTB_INDEX3_LO          : 9'h012        ,
	BTB_SIZE               : 14'h0200      ,
	BTB_TOFFSET_SIZE       : 9'h00C        ,
	BUILD_AHB_LITE         : 4'h0          ,
	BUILD_AXI4             : 5'h01         ,
	BUILD_AXI_NATIVE       : 5'h01         ,
	BUS_PRTY_DEFAULT       : 6'h03         ,
	DATA_ACCESS_ADDR0      : 36'h000000000  ,
	DATA_ACCESS_ADDR1      : 36'h000000000  ,
	DATA_ACCESS_ADDR2      : 36'h000000000  ,
	DATA_ACCESS_ADDR3      : 36'h000000000  ,
	DATA_ACCESS_ADDR4      : 36'h000000000  ,
	DATA_ACCESS_ADDR5      : 36'h000000000  ,
	DATA_ACCESS_ADDR6      : 36'h000000000  ,
	DATA_ACCESS_ADDR7      : 36'h000000000  ,
	DATA_ACCESS_ENABLE0    : 5'h00         ,
	DATA_ACCESS_ENABLE1    : 5'h00         ,
	DATA_ACCESS_ENABLE2    : 5'h00         ,
	DATA_ACCESS_ENABLE3    : 5'h00         ,
	DATA_ACCESS_ENABLE4    : 5'h00         ,
	DATA_ACCESS_ENABLE5    : 5'h00         ,
	DATA_ACCESS_ENABLE6    : 5'h00         ,
	DATA_ACCESS_ENABLE7    : 5'h00         ,
	DATA_ACCESS_MASK0      : 36'h0FFFFFFFF  ,
	DATA_ACCESS_MASK1      : 36'h0FFFFFFFF  ,
	DATA_ACCESS_MASK2      : 36'h0FFFFFFFF  ,
	DATA_ACCESS_MASK3      : 36'h0FFFFFFFF  ,
	DATA_ACCESS_MASK4      : 36'h0FFFFFFFF  ,
	DATA_ACCESS_MASK5      : 36'h0FFFFFFFF  ,
	DATA_ACCESS_MASK6      : 36'h0FFFFFFFF  ,
	DATA_ACCESS_MASK7      : 36'h0FFFFFFFF  ,
	DCCM_BANK_BITS         : 7'h02         ,
	DCCM_BITS              : 9'h010        ,
	DCCM_BYTE_WIDTH        : 7'h04         ,
	DCCM_DATA_WIDTH        : 10'h020        ,
	DCCM_ECC_WIDTH         : 7'h07         ,
	DCCM_ENABLE            : 5'h01         ,
	DCCM_FDATA_WIDTH       : 10'h027        ,
	DCCM_INDEX_BITS        : 8'h0C         ,
	DCCM_NUM_BANKS         : 9'h004        ,
	DCCM_REGION            : 8'h0F         ,
	DCCM_SADR              : 36'h0F0040000  ,
	DCCM_SIZE              : 14'h0040       ,
	DCCM_WIDTH_BITS        : 6'h02         ,
	DIV_BIT                : 7'h04         ,
	DIV_NEW                : 5'h01         ,
	DMA_BUF_DEPTH          : 7'h05         ,
	DMA_BUS_ID             : 9'h001        ,
	DMA_BUS_PRTY           : 6'h02         ,
	DMA_BUS_TAG            : 8'h01         ,
	FAST_INTERRUPT_REDIRECT : 5'h01         ,
	ICACHE_2BANKS          : 5'h01         ,
	ICACHE_BANK_BITS       : 7'h01         ,
	ICACHE_BANK_HI         : 7'h03         ,
	ICACHE_BANK_LO         : 6'h03         ,
	ICACHE_BANK_WIDTH      : 8'h08         ,
	ICACHE_BANKS_WAY       : 7'h02         ,
	ICACHE_BEAT_ADDR_HI    : 8'h05         ,
	ICACHE_BEAT_BITS       : 8'h03         ,
	ICACHE_BYPASS_ENABLE   : 5'h01         ,
	ICACHE_DATA_DEPTH      : 18'h00200      ,
	ICACHE_DATA_INDEX_LO   : 7'h04         ,
	ICACHE_DATA_WIDTH      : 11'h040        ,
	ICACHE_ECC             : 5'h01         ,
	ICACHE_ENABLE          : 5'h01         ,
	ICACHE_FDATA_WIDTH     : 11'h047        ,
	ICACHE_INDEX_HI        : 9'h00C        ,
	ICACHE_LN_SZ           : 11'h040        ,
	ICACHE_NUM_BEATS       : 8'h08         ,
	ICACHE_NUM_BYPASS      : 8'h02         ,
	ICACHE_NUM_BYPASS_WIDTH : 8'h02         ,
	ICACHE_NUM_WAYS        : 7'h02         ,
	ICACHE_ONLY            : 5'h00         ,
	ICACHE_SCND_LAST       : 8'h06         ,
	ICACHE_SIZE            : 13'h0010       ,
	ICACHE_STATUS_BITS     : 7'h01         ,
	ICACHE_TAG_BYPASS_ENABLE : 5'h01         ,
	ICACHE_TAG_DEPTH       : 17'h00080      ,
	ICACHE_TAG_INDEX_LO    : 7'h06         ,
	ICACHE_TAG_LO          : 9'h00D        ,
	ICACHE_TAG_NUM_BYPASS  : 8'h02         ,
	ICACHE_TAG_NUM_BYPASS_WIDTH : 8'h02         ,
	ICACHE_WAYPACK         : 5'h01         ,
	ICCM_BANK_BITS         : 7'h02         ,
	ICCM_BANK_HI           : 9'h003        ,
	ICCM_BANK_INDEX_LO     : 9'h004        ,
	ICCM_BITS              : 9'h010        ,
	ICCM_ENABLE            : 5'h01         ,
	ICCM_ICACHE            : 5'h01         ,
	ICCM_INDEX_BITS        : 8'h0C         ,
	ICCM_NUM_BANKS         : 9'h004        ,
	ICCM_ONLY              : 5'h00         ,
	ICCM_REGION            : 8'h0E         ,
	ICCM_SADR              : 36'h0EE000000  ,
	ICCM_SIZE              : 14'h0040       ,
	IFU_BUS_ID             : 5'h01         ,
	IFU_BUS_PRTY           : 6'h02         ,
	IFU_BUS_TAG            : 8'h03         ,
	INST_ACCESS_ADDR0      : 36'h000000000  ,
	INST_ACCESS_ADDR1      : 36'h000000000  ,
	INST_ACCESS_ADDR2      : 36'h000000000  ,
	INST_ACCESS_ADDR3      : 36'h000000000  ,
	INST_ACCESS_ADDR4      : 36'h000000000  ,
	INST_ACCESS_ADDR5      : 36'h000000000  ,
	INST_ACCESS_ADDR6      : 36'h000000000  ,
	INST_ACCESS_ADDR7      : 36'h000000000  ,
	INST_ACCESS_ENABLE0    : 5'h00         ,
	INST_ACCESS_ENABLE1    : 5'h00         ,
	INST_ACCESS_ENABLE2    : 5'h00         ,
	INST_ACCESS_ENABLE3    : 5'h00         ,
	INST_ACCESS_ENABLE4    : 5'h00         ,
	INST_ACCESS_ENABLE5    : 5'h00         ,
	INST_ACCESS_ENABLE6    : 5'h00         ,
	INST_ACCESS_ENABLE7    : 5'h00         ,
	INST_ACCESS_MASK0      : 36'h0FFFFFFFF  ,
	INST_ACCESS_MASK1      : 36'h0FFFFFFFF  ,
	INST_ACCESS_MASK2      : 36'h0FFFFFFFF  ,
	INST_ACCESS_MASK3      : 36'h0FFFFFFFF  ,
	INST_ACCESS_MASK4      : 36'h0FFFFFFFF  ,
	INST_ACCESS_MASK5      : 36'h0FFFFFFFF  ,
	INST_ACCESS_MASK6      : 36'h0FFFFFFFF  ,
	INST_ACCESS_MASK7      : 36'h0FFFFFFFF  ,
	LOAD_TO_USE_PLUS1      : 5'h00         ,
	LSU2DMA                : 5'h00         ,
	LSU_BUS_ID             : 5'h01         ,
	LSU_BUS_PRTY           : 6'h02         ,
	LSU_BUS_TAG            : 8'h03         ,
	LSU_NUM_NBLOAD         : 9'h004        ,
	LSU_NUM_NBLOAD_WIDTH   : 7'h02         ,
	LSU_SB_BITS            : 9'h010        ,
	LSU_STBUF_DEPTH        : 8'h04         ,
	NO_ICCM_NO_ICACHE      : 5'h00         ,
	PIC_2CYCLE             : 5'h00         ,
	PIC_BASE_ADDR          : 36'h0F00C0000  ,
	PIC_BITS               : 9'h00F        ,
	PIC_INT_WORDS          : 8'h01         ,
	PIC_REGION             : 8'h0F         ,
	PIC_SIZE               : 13'h0020       ,
	PIC_TOTAL_INT          : 12'h01F        ,
	PIC_TOTAL_INT_PLUS1    : 13'h0020       ,
	RET_STACK_SIZE         : 8'h08         ,
	SB_BUS_ID              : 5'h01         ,
	SB_BUS_PRTY            : 6'h02         ,
	SB_BUS_TAG             : 8'h01         ,
	TIMER_LEGAL_EN         : 5'h01         
}
