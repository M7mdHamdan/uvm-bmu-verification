typedef enum {Actual, Expected} itemKind;